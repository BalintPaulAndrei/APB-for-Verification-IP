package rst_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"
    `include "rst_item.svh"
    `include "rst_monitor.svh"
    `include "rst_driver.svh"
    `include "rst_sequencer.svh"
    `include "rst_agent.svh"
    `include "rst_sequence.svh"

endpackage : rst_pkg