package afvip_tb_pkg;
            
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import apb_pkg::*;
    import intr_pkg::*;
    import rst_pkg::*;

   
    `include "afvip_scoreboard.svh"
    `include "afvip_coverage.svh"
    `include "afvip_environment.svh"

endpackage : afvip_tb_pkg