// -----------------------------------------------------------------------------
// Module name: rst_if
// HDL        : System Verilog
// Author     : Balint Paul
// Description: Encapsulate signals into a block
// Date       : 28 June 2023
// -----------------------------------------------------------------------------
interface rst_if(
    input     clk,       // clk
    input reg reset      // reset
)
    
    import uvm_pkg::*;
    //logic reset;
    

endinterface : rst_if