package afvip_test_pkg;

    import uvm_pkg::*;
    import apb_pkg::*;
    import intr_pkg::*;
    import rst_pkg::*;
    import afvip_tb_pkg::*;
    
    `include "uvm_macros.svh"
    `include "afvip_test_lib.svh"

endpackage : afvip_test_pkg