package intr_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"
    `include "intr_item.svh"
    `include "intr_monitor.svh"
    `include "intr_agent.svh"

endpackage : intr_pkg